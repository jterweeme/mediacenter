module va1(
    input csi_clk,
    input csi_reset_n,
    
    output wire avs_s1_

