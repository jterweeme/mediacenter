module myvgascratch1(
    input csi_clk_sys,
    input csi_reset_n,
    input csi_clk25);

always @

endmodule


