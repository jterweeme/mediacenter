module toetsenbord2(
    clk
);


