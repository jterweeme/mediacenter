LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_misc.all;

-- ******************************************************************************
-- * License Agreement                                                          *
-- *                                                                            *
-- * Copyright (c) 1991-2013 Altera Corporation, San Jose, California, USA.     *
-- * All rights reserved.                                                       *
-- *                                                                            *
-- * Any megafunction design, and related net list (encrypted or decrypted),    *
-- *  support information, device programming or simulation file, and any other *
-- *  associated documentation or information provided by Altera or a partner   *
-- *  under Altera's Megafunction Partnership Program may be used only to       *
-- *  program PLD devices (but not masked PLD devices) from Altera.  Any other  *
-- *  use of such megafunction design, net list, support information, device    *
-- *  programming or simulation file, or any other related documentation or     *
-- *  information is prohibited for any other purpose, including, but not       *
-- *  limited to modification, reverse engineering, de-compiling, or use with   *
-- *  any other silicon devices, unless such use is explicitly licensed under   *
-- *  a separate agreement with Altera or a megafunction partner.  Title to     *
-- *  the intellectual property, including patents, copyrights, trademarks,     *
-- *  trade secrets, or maskworks, embodied in any such megafunction design,    *
-- *  net list, support information, device programming or simulation file, or  *
-- *  any other related documentation or information provided by Altera or a    *
-- *  megafunction partner, remains with Altera, the megafunction partner, or   *
-- *  their respective licensors.  No other licenses, including any licenses    *
-- *  needed under any third party's intellectual property, are provided herein.*
-- *  Copying or modifying any file, or portion thereof, to which this notice   *
-- *  is attached violates this copyright.                                      *
-- *                                                                            *
-- * THIS FILE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR    *
-- * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,   *
-- * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL    *
-- * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER *
-- * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING    *
-- * FROM, OUT OF OR IN CONNECTION WITH THIS FILE OR THE USE OR OTHER DEALINGS  *
-- * IN THIS FILE.                                                              *
-- *                                                                            *
-- * This agreement shall be governed in all respects by the laws of the State  *
-- *  of California and by the laws of the United States of America.            *
-- *                                                                            *
-- ******************************************************************************

-- ******************************************************************************
-- *                                                                            *
-- * This module reads and writes data to USB chip on the DE2 Board.            *
-- *                                                                            *
-- ******************************************************************************

ENTITY Altera_UP_Avalon_USB IS 

-- *****************************************************************************
-- *                             Generic Declarations                          *
-- *****************************************************************************

-- *****************************************************************************
-- *                             Port Declarations                             *
-- *****************************************************************************
PORT (
	-- Inputs
	clk				:IN		STD_LOGIC;
	reset				:IN		STD_LOGIC;

	address			:IN		STD_LOGIC_VECTOR( 1 DOWNTO  0);	
	chipselect		:IN		STD_LOGIC;
	read				:IN		STD_LOGIC;
	write				:IN		STD_LOGIC;
	writedata		:IN		STD_LOGIC_VECTOR(15 DOWNTO  0);	

	OTG_INT0			:IN		STD_LOGIC;
	OTG_INT1			:IN		STD_LOGIC;

	-- Bidirectionals
	OTG_DATA			:INOUT	STD_LOGIC_VECTOR(15 DOWNTO  0);	

	-- Outputs
	readdata			:BUFFER	STD_LOGIC_VECTOR(15 DOWNTO  0);	

	irq				:BUFFER	STD_LOGIC;

	OTG_RST_N		:BUFFER	STD_LOGIC;
	OTG_ADDR			:BUFFER	STD_LOGIC_VECTOR( 1 DOWNTO  0);	
	OTG_CS_N			:BUFFER	STD_LOGIC;
	OTG_RD_N			:BUFFER	STD_LOGIC;
	OTG_WR_N			:BUFFER	STD_LOGIC

);

END Altera_UP_Avalon_USB;

ARCHITECTURE Behaviour OF Altera_UP_Avalon_USB IS
-- *****************************************************************************
-- *                           Constant Declarations                           *
-- *****************************************************************************

-- *****************************************************************************
-- *                       Internal Signals Declarations                       *
-- *****************************************************************************
	-- Internal Wires
	
	-- Internal Registers
	SIGNAL	data_to_usb_chip	:STD_LOGIC_VECTOR(15 DOWNTO  0);	
	
	-- State Machine Registers
	
-- *****************************************************************************
-- *                          Component Declarations                           *
-- *****************************************************************************
BEGIN
-- *****************************************************************************
-- *                         Finite State Machine(s)                           *
-- *****************************************************************************


-- *****************************************************************************
-- *                             Sequential Logic                              *
-- *****************************************************************************

	PROCESS (clk)
	BEGIN
		IF clk'EVENT AND clk = '1' THEN
			IF (reset = '1') THEN
				readdata				<= B"0000000000000000";
		
				irq					<= '0';
		
				data_to_usb_chip	<= B"0000000000000000";
		
				OTG_RST_N			<= '0';
				OTG_ADDR				<= B"00";
				OTG_CS_N				<= '1';
				OTG_RD_N				<= '1';
				OTG_WR_N				<= '1';
			ELSE
				readdata				<= OTG_DATA;
		
				irq					<= NOT OTG_INT1 OR NOT OTG_INT0;
				
				data_to_usb_chip	<= writedata(15 DOWNTO 0);
		
				OTG_RST_N			<= '1';
				OTG_ADDR				<= address;
				OTG_CS_N				<= NOT chipselect;
				OTG_RD_N				<= NOT read;
				OTG_WR_N				<= NOT write;
			END IF;
		END IF;
	END PROCESS;


-- *****************************************************************************
-- *                            Combinational Logic                            *
-- *****************************************************************************

	OTG_DATA <= (OTHERS => 'Z') WHEN (OTG_WR_N = '1') ELSE data_to_usb_chip;

-- *****************************************************************************
-- *                          Component Instantiations                         *
-- *****************************************************************************



END Behaviour;
