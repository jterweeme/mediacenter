module myi2c1(
    
);
