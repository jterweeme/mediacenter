module infrared(iCLK, iRST_n, iIRDA, iREAD,
                    oDATA_REAY,
                    oDATA);

input iCLK, iRST_n, iIRDA, iREAD, oDATA_REAY, oDATA;
                    
endmodule

